class aux_seqr extends uvm_sequencer#(aux_xtn);
`uvm_component_utils(aux_seqr);
function new(string name="aux_seqr",uvm_component parent);
super.new(name,parent);
endfunction
endclass
